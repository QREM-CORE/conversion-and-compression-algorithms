module tb_byte_encode;
endmodule