module tb_bytes2bits;
endmodule