module byte_decode;
endmodule