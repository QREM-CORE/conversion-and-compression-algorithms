module tb_byte_decode;
endmodule