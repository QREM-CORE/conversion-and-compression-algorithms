module bits2bytes;
endmodule