module byte_encode;
endmodule