module tb_bits2bytes;
endmodule