module bytes2bits;
endmodule